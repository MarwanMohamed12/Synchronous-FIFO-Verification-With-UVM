package shared_pkg;
    int error_count, correct_count;   
endpackage


